package TagEngine(MkTagType) where

type MkTagType inFlightTransactions = UInt (TLog inFlightTransactions)
