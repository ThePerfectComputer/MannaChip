package TransactionToSubtransaction(
    Len, Offset, DeviceLine,
    Subtransaction(..),
    TransactionToSubtransactionAdapter(..),
    mkTransactionToSubtransactionAdapter) where

import SpecialFIFOs
import FIFO
import Words
import BusTypes
import TagEngine

type Len        = UInt 5 -- a subtransaction can be up to 16 bytes long in length
type Offset     = UInt 4 -- and can be offset by up to 15 bytes
type DeviceLine = Addr   -- address of device line for given subtransaction

data Subtransaction = NonTerminating    DeviceLine Offset Len
                    | Terminating       DeviceLine Offset Len
                    deriving (Bits, FShow, Eq)

subtransactionLen :: Subtransaction -> Len
subtransactionLen (NonTerminating _ _ len) = len
subtransactionLen (Terminating    _ _ len) = len

nextSubtransaction :: Addr -> Addr -> (Maybe Addr) -> WordSize -> Subtransaction
nextSubtransaction startAddr endAddr previousAddr deviceLineSize =
    let
        shiftAmt :: Integer
        shiftAmt = wordSizeToAddrShiftAmt deviceLineSize

        currAddr :: Addr
        currAddr = case previousAddr of
            Just addr -> addr
            Nothing -> startAddr

        currLineAddrDeviceSpace :: DeviceLine
        currLineAddrDeviceSpace = currAddr >> shiftAmt

        lineAddrLeftBoundBusSpace :: Addr
        lineAddrLeftBoundBusSpace = currLineAddrDeviceSpace << shiftAmt

        lineAddrRightBoundBusSpace :: Addr
        lineAddrRightBoundBusSpace = (currLineAddrDeviceSpace + 1) << shiftAmt

        offset :: Offset
        offset = truncate $ currAddr - lineAddrLeftBoundBusSpace

        len :: Len
        len = truncate $
            min (endAddr - currAddr) (lineAddrRightBoundBusSpace - currAddr)

        terminating :: Bool
        terminating = endAddr == currAddr + (zeroExtend len)
    in
        case terminating of
            True  -> Terminating currLineAddrDeviceSpace offset len
            False -> NonTerminating currLineAddrDeviceSpace offset len

transactionRequestToAddr :: TransactionRequest -> Addr
transactionRequestToAddr (ReadRequest addr _) = addr
transactionRequestToAddr (WriteRequest addr _) = addr

transactionDataToWordSize :: TransactionData -> WordSize
transactionDataToWordSize (Byte _)          = Words.Byte
transactionDataToWordSize (HalfWord _)      = Words.HalfWord
transactionDataToWordSize (FullWord _)      = Words.FullWord
transactionDataToWordSize (DoubleWord _)    = Words.DoubleWord
transactionDataToWordSize (QuadWord _)      = Words.QuadWord

transactionRequestToWordSize :: TransactionRequest -> WordSize
transactionRequestToWordSize (ReadRequest  _ s) = s
transactionRequestToWordSize (WriteRequest _ d) = transactionDataToWordSize d

interface (TransactionToSubtransactionAdapter:: # -> *) inFlightTransactions =
    {
    enqueueTransaction      :: (TaggedTransactionRequest inFlightTransactions) -> Action;
    dequeueSubTransaction   :: ActionValue Subtransaction;
    currentTransactionTag   :: MkTagType inFlightTransactions;
    }

mkTransactionToSubtransactionAdapter ::
    WordSize ->
    Module (TransactionToSubtransactionAdapter inFlightTransactions)
mkTransactionToSubtransactionAdapter deviceLineSize = do

    transactionQueue :: FIFO (TaggedTransactionRequest inFlightTransactions)
    transactionQueue <- mkBypassFIFO

    subTransactionQueue :: FIFO Subtransaction
    subTransactionQueue <- mkBypassFIFO

    previousAddr :: Reg (Maybe Addr)
    previousAddr <- mkReg Nothing

    let startAddr :: Addr
        startAddr =  transactionRequestToAddr $ transactionQueue.first.request

        endAddr :: Addr
        endAddr = startAddr + (
            fromInteger $ wordSizeNumBytes $
            transactionRequestToWordSize transactionQueue.first.request
            )

    addRules $
      rules
        "nextSubtransaction" : when True ==>
            do
                let
                    subtransaction :: Subtransaction
                    subtransaction =
                        nextSubtransaction startAddr endAddr previousAddr deviceLineSize

                    subtransactionLenVal :: Addr
                    subtransactionLenVal = zeroExtend $ subtransactionLen subtransaction

                subTransactionQueue.enq subtransaction

                case subtransaction of
                    NonTerminating _ _ _ ->
                        do
                            previousAddr := case previousAddr of
                                Just addr -> Just $ addr + subtransactionLenVal
                                Nothing   -> Just $ startAddr + subtransactionLenVal
                    Terminating _ _ _ ->
                        do
                            previousAddr := Nothing
                            transactionQueue.deq

    return $
        interface TransactionToSubtransactionAdapter
            enqueueTransaction  :: (TaggedTransactionRequest inFlightTransactions) -> Action
            enqueueTransaction taggedTransactionRequest =
                transactionQueue.enq taggedTransactionRequest

            dequeueSubTransaction   :: ActionValue Subtransaction
            dequeueSubTransaction = do
                subTransactionQueue.deq
                return subTransactionQueue.first

            currentTransactionTag   :: MkTagType inFlightTransactions
            currentTransactionTag = transactionQueue.first.tag
