package Top(mkTop, ITop(..)) where

import Deserializer
import Core
import Serializer
import BRAM
import CBindings

type FCLK = 25000000
type BAUD = 9600

interface ITop = {
  ftdi_rxd :: Bit 1           {-# always_ready  #-}
 ;led      :: Bit 8           {-# always_ready  #-}
 ;ftdi_txd :: Bit 1 -> Action {-# always_ready , always_enabled  #-}
};

mkTop :: Module ITop
mkTop = do
  fileHandle   :: Handle <- openFile "compile.log" WriteMode
  deserializer :: IDeserializer FCLK BAUD <- mkDeserialize fileHandle
  serializer   :: ISerializer FCLK BAUD <- mkSerialize fileHandle
  core         :: Core FCLK <- mkCore
  persistLed  :: Reg (Bit 8) <- mkReg 0
  messageM $ "Hallo!!" + (realToString 5)

  -- refactor such that the following rules are let-bound to 
  -- `attachIO` identifier
  addRules $
    rules
      "coreLedO" : when True ==>
        persistLed := core.getLed

      "coreCharDeviceO" : when True ==>
        serializer.putBit8 core.getChar

      "coreCharDeviceO" : when True ==>
        serializer.putBit8 core.getChar

      "coreCharDeviceI" : when True ==>
        core.putChar deserializer.get

  return $
    interface ITop
      ftdi_rxd =  serializer.bitLineOut
      ftdi_txd bitIn =  
           do
             deserializer.putBitIn bitIn
      led =  persistLed

mkSim :: Module Empty
mkSim = do
  let cfg          :: BRAM_Configure = defaultValue

  count            :: Reg (UInt 3) <- mkReg 0;
  initCFunctions :: Reg Bool <- mkReg False;
  core             :: Core FCLK <- mkCore;

  addRules $
    rules
      "initCFunctionsOnce":  when not initCFunctions ==>
        do
          initTerminal
          setupSigintHandler
          initCFunctions := True
      "coreCharDeviceO":  when True ==>
        do
          writeCharToTerminal core.getChar
      "coreCharDeviceI":  when (isCharAvailable == 1) ==>
        do
          core.putChar getCharFromTerminal
      "endSim":  when wasCtrlCReceived ==>
        do
          restoreTerminal
          $display "GOT CTRL+C"
          $finish