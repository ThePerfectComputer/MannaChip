package Top(mkTop, ITop(..)) where

import Deserializer
import Serializer
import CBindings
import BusTypes

type UART_CLK_PERIOD = 2604 -- for 9600 BAUD at 25MHz

interface ITop = {
  ftdi_rxd :: Bit 1           {-# always_ready  #-}
 ;led      :: Bit 8           {-# always_ready  #-}
 ;ftdi_txd :: Bit 1 -> Action {-# always_ready , always_enabled  #-}
};

mkTop :: Module ITop
mkTop = do
  fileHandle   :: Handle <- openFile "compile.log" WriteMode
  deserializer :: IDeserializer UART_CLK_PERIOD <- mkDeserialize fileHandle
  serializer   :: ISerializer UART_CLK_PERIOD <- mkSerialize fileHandle
  recentByte   :: Reg (Bit 8) <- mkReg 0
  messageM $ "Hallo!!" + (realToString 5)

  addRules $
    rules
      "loopback" : when True ==>
        do
          let byte = deserializer.get
          recentByte := byte
          serializer.putBit8 byte

  return $
    interface ITop
      ftdi_rxd =  serializer.bitLineOut
      ftdi_txd bitIn =
           do
             deserializer.putBitIn bitIn
      led =  recentByte

mkSim :: Module Empty
mkSim = do
  initCFunctions :: Reg Bool <- mkReg False;

  addRules $
    rules
      "initCFunctionsOnce":  when not initCFunctions ==>
        do
          initTerminal
          setupSigintHandler
          initCFunctions := True

      "loopback":  when (isCharAvailable == 1) ==>
        do
          writeCharToTerminal getCharFromTerminal

      "endSim":  when wasCtrlCReceived ==>
        do
          restoreTerminal
          $display "GOT CTRL+C"
          $finish
