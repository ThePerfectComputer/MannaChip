package BusTypes(
    Addr,
    BusError(..),
    TransactionData(..),
    TransactionRequest(..),
    TransactionResponse(..),
    TaggedTransactionRequest(..),
    TaggedTransactionResponse(..)) where

import TagEngine
import Words

type Addr = UInt 64

data BusError = MisAligned Addr
                deriving (Bits, FShow, Eq)

data TransactionData = Byte (UInt 8)
                     | HalfWord (UInt 16)
                     | FullWord (UInt 32)
                     | DoubleWord (UInt 64)
                     | QuadWord (UInt 128)
                     deriving (Bits, FShow, Eq)

data TransactionRequest = ReadRequest  Addr WordSize
                        | WriteRequest Addr TransactionData
                        deriving (Bits, FShow, Eq)

data TransactionResponse = ReadResponse  (Either BusError TransactionData)
                         | WriteResponse (Either BusError ())
                         deriving (Bits, FShow, Eq)


struct TaggedTransactionRequest inFlightTransactions =
    { tag       :: MkTagType inFlightTransactions;
      request   :: TransactionRequest
    }
    deriving (Bits, FShow, Eq)

struct TaggedTransactionResponse inFlightTransactions =
    { tag       :: MkTagType inFlightTransactions;
      response  :: TransactionResponse
    }
    deriving (Bits, FShow, Eq)
